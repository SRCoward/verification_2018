module sam_log2(X,k,z);
parameter y_width=6;
input [22:0] X;
input [5:0] k;
output [22:0] z;
wire [5:0] y;
wire [17:0] x;
reg [13:0] a;
reg [37:0] b;
reg [60:0] c;
wire [34:0] x_hat;
wire [120:0] t;
wire [120:0] s;
wire [120:0] zz;
assign k=0;
assign y=X[22:17];
assign x=X[16:0];

always @ (y) begin
	case(y)
		6'B000000:begin a=14'B10110101110101; b=38'B10111000101010000101011101000010101110; c=60'B0; end
		6'B000001:begin a=14'B10110000010100; b=38'B10110101110100010010000101100011011000; c=60'B1011011100111100101101000010111000010110100100010101000; end
		6'B000010:begin a=14'B10101011000011; b=38'B10110011000011111111010001000101001111; c=60'B10110101110101101001101110101100011101111110110000111000; end
		6'B000011:begin a=14'B10100110000001; b=38'B10110000011000111101001101011111011111; c=60'B100001110101100111000100111111010001010011111100110110000; end
		6'B000100:begin a=14'B10100001001110; b=38'B10101101110010111101000100000011100011; c=60'B101100110001111110110111110101100100100010011000101100000; end
		6'B000101:begin a=14'B10011100100111; b=38'B10101011010001110000110101001001100100; c=60'B110111100100001000010010000001010110110101011101110110000; end
		6'B000110:begin a=14'B10011000001100; b=38'B10101000110101001011010100010100100100; c=60'B1000010001100010110001000110011011010011110011110010000000; end
		6'B000111:begin a=14'B10010011111110; b=38'B10100110011101000000000100101011110111; c=60'B1001100101010111010011110001001111000101011100001101000000; end
		6'B001000:begin a=14'B10001111111010; b=38'B10100100001001000011010101100111101100; c=60'B1010111000000000110100011100111111011110101101000100000000; end
		6'B001001:begin a=14'B10001100000010; b=38'B10100001111001001001111111101111001101; c=60'B1100001001100001010111101000000101111000000111011001100000; end
		6'B001010:begin a=14'B10001000010011; b=38'B10011111101101001001100010000110001111; c=60'B1101011001111010111100010110110110100111011001001010000000; end
		6'B001011:begin a=14'B10000100101101; b=38'B10011101100100110111111111101001001110; c=60'B1110101001001111011100100110000110010010110010110111100000; end
		6'B001100:begin a=14'B10000001010001; b=38'B10011011100000001011111100110110001010; c=60'B1111110111100000101101011100100000010011010000000101100000; end
		6'B001101:begin a=14'B1111101111100; b=38'B10011001011110111100011101100001011000; c=60'B10001000100110000011111011010110100110000101101110110000000; end
		6'B001110:begin a=14'B1111010110000; b=38'B10010111100001000001000010110100110011; c=60'B10010010001000000011110101011000011100000011100111001000000; end
		6'B001111:begin a=14'B1110111101100; b=38'B10010101100110010001101001011001010001; c=60'B10011011100010010010011001110101001001100110111101101000000; end
		6'B010000:begin a=14'B1110100101111; b=38'B10010011101110100110100111101000100011; c=60'B10100100110100111100001001011110011010001101110001011000000; end
		6'B010001:begin a=14'B1110001111001; b=38'B10010001111001111000101100000111100111; c=60'B10101110000000001101000111001111110111101011010001000000000; end
		6'B010010:begin a=14'B1101111001001; b=38'B10010000001000000000111100001000001110; c=60'B10110111000100010000111001101100111010000110011011111000000; end
		6'B010011:begin a=14'B1101100100000; b=38'B10001110011000111000110010010001100010; c=60'B11000000000001010010101100011000101100001110001010100000000; end
		6'B010100:begin a=14'B1101001111100; b=38'B10001100101100011001111101001110110010; c=60'B11001000110111011101010001001000111110001011100001001000000; end
		6'B010101:begin a=14'B1100111011111; b=38'B10001011000010011110011110100011101110; c=60'B11010001100110111011000001010011111110110000001010001000000; end
		6'B010110:begin a=14'B1100101000110; b=38'B10001001011011000000101001100110011101; c=60'B11011010001111110101111110111001110001000001010100001000000; end
		6'B010111:begin a=14'B1100010110011; b=38'B10000111110101111011000010011101111100; c=60'B11100010110010010111110101101001010010101101101010111000000; end
		6'B011000:begin a=14'B1100000100101; b=38'B10000110010011001000011101000101000111; c=60'B11101011001110101001111100000001100101110101000001111000000; end
		6'B011001:begin a=14'B1011110011100; b=38'B10000100110010100011111100010001111101; c=60'B11110011100100110101010100001111001110101010011010010000000; end
		6'B011010:begin a=14'B1011100010111; b=38'B10000011010100001000110001000000100010; c=60'B11111011110101000010101101000110010110000011011001111000000; end
		6'B011011:begin a=14'B1011010010111; b=38'B10000001110111110010011001100001011000; c=60'B100000011111111011010100010111001011110011001100000000000000; end
		6'B011100:begin a=14'B1011000011010; b=38'B10000000011101011100100000101011001100; c=60'B100001100000100000101000000001101011000111010101001110000000; end
		6'B011101:begin a=14'B1010110100010; b=38'B1111111000101000010111101001111011110; c=60'B100010100000011001001111110101010000111100101010000110000000; end
		6'B011110:begin a=14'B1010100101101; b=38'B1111101101110100001110001010010000001; c=60'B100011011111100110001000111101001010111010000000011100000000; end
		6'B011111:begin a=14'B1010010111100; b=38'B1111100011001110101001001100010110100; c=60'B100100011110001000001110101000010011100100111110010000000000; end
		6'B100000:begin a=14'B1010001001111; b=38'B1111011000110111001011100111010011111; c=60'B100101011100000000011010001110011111101111010110100010000000; end
		6'B100001:begin a=14'B1001111100101; b=38'B1111001110101101011001011111000110110; c=60'B100110011001001111100011010101011010010011100101001110000000; end
		6'B100010:begin a=14'B1001101111110; b=38'B1111000100110000111000000000101011110; c=60'B100111010101110110011111110101010000000100001011001110000000; end
		6'B100011:begin a=14'B1001100011010; b=38'B1110111011000001001101011110010010001; c=60'B101000010001110110000011111101001100001101010101010100000000; end
		6'B100100:begin a=14'B1001010111001; b=38'B1110110001011110000001001011111101111; c=60'B101001001101001111000010010111100110100011011100010110000000; end
		6'B100101:begin a=14'B1001001011011; b=38'B1110101000000110111011011100010111100; c=60'B101010001000000010001100001110000100010101000111110010000000; end
		6'B100110:begin a=14'B1001000000000; b=38'B1110011110111011100101011101100111001; c=60'B101011000010010000010001001101001100010011101001101000000000; end
		6'B100111:begin a=14'B1000110101000; b=38'B1110010101111011101001010110011100011; c=60'B101011111011111001111111101000001111000001001101011110000000; end
		6'B101000:begin a=14'B1000101010001; b=38'B1110001101000110110010000011011111110; c=60'B101100110101000000000100011100100011110001000110011000000000; end
		6'B101001:begin a=14'B1000011111110; b=38'B1110000100011100101011010100101110011; c=60'B101101101101100011001011010100111011000011001010010100000000; end
		6'B101010:begin a=14'B1000010101101; b=38'B1101111011111101000001101010111111010; c=60'B101110100101100011111110101100100111000000111010101000000000; end
		6'B101011:begin a=14'B1000001011110; b=38'B1101110011100111100010010101110001010; c=60'B101111011101000011000111110010011010100000010111001000000000; end
		6'B101100:begin a=14'B1000000010001; b=38'B1101101011011011111011010001000000100; c=60'B110000010100000001001110101011011111001110000011100110000000; end
		6'B101101:begin a=14'B111111000110; b=38'B1101100011011001111011000011000011111; c=60'B110001001010011110111010010110000011011101111100010110000000; end
		6'B101110:begin a=14'B111101111101; b=38'B1101011011100001010000111010110010011; c=60'B110010000000011100110000101100000000000000010110011100000000; end
		6'B101111:begin a=14'B111100110110; b=38'B1101010011110001101100101101101101010; c=60'B110010110101111011010110100101010110010110101111101100000000; end
		6'B110000:begin a=14'B111011110001; b=38'B1101001100001010111110110110010010101; c=60'B110011101010111011001111111010101000000010000101100110000000; end
		6'B110001:begin a=14'B111010101110; b=38'B1101000100101100111000010010010011111; c=60'B110100011111011100111111100111000111000011000001000000000000; end
		6'B110010:begin a=14'B111001101101; b=38'B1100111101010111001010100001010011011; c=60'B110101010011100001000111101011000000000010100110101000000000; end
		6'B110011:begin a=14'B111000101101; b=38'B1100110110001001100111100011000110010; c=60'B110110000111001000001001001101011110011001000011011000000000; end
		6'B110100:begin a=14'B110111101111; b=38'B1100101111000100000001110110011011000; c=60'B110110111010010010100100011110101010100110010110110100000000; end
		6'B110101:begin a=14'B110110110011; b=38'B1100101000000110001100010111100101010; c=60'B110111101101000000111000111001100011001111110011011100000000; end
		6'B110110:begin a=14'B110101111000; b=38'B1100100001001111111010011111001110000; c=60'B111000011111010011100101000101110000110100000010101100000000; end
		6'B110111:begin a=14'B110100111110; b=38'B1100011010100001000000000001000110011; c=60'B111001010001001011000110111001010100100110011000101110000000; end
		6'B111000:begin a=14'B110100000110; b=38'B1100010011111001010001001011000000011; c=60'B111010000010100111111011011010010011000001000100101100000000; end
		6'B111001:begin a=14'B110011010000; b=38'B1100001101011000100010100011101001011; c=60'B111010110011101010011111000000011001011101010000011110000000; end
		6'B111010:begin a=14'B110010011010; b=38'B1100000110111110101001001001101001000; c=60'B111011100100010011001101010110011111111110101011011010000000; end
		6'B111011:begin a=14'B110001100110; b=38'B1100000000101011011010010010100011000; c=60'B111100010100100010100001011100000111000000001010000010000000; end
		6'B111100:begin a=14'B110000110100; b=38'B1011111010011110101011101001111011111; c=60'B111101000100011000110101100110110001001101010011100110000000; end
		6'B111101:begin a=14'B110000000010; b=38'B1011110100011000010011010000100000101; c=60'B111101110011110110100011100011011001110101001010100000000000; end
		6'B111110:begin a=14'B101111010010; b=38'B1011101110011000000111011011010001010; c=60'B111110100010111100000100010111100111100000110010101100000000; end
		6'B111111:begin a=14'B101110100010; b=38'B1011101000011101111110110010101101000; c=60'B111111010001101001110000100010111011111000010001100110000000; end
	endcase
end
assign x_hat=(x*x)<<60;
assign t=a*(x_hat>>k);
assign s = b*(x<<60);
//assign t=(x*x)>>k;
assign zz=s-t+(c<<60);
	
assign z=(zz>>97);

endmodule
